module module_name(
    sys_clk    ,
    sys_rst_n  ,
    
);

input               sys_clk;
input               sys_rst_n;


endmodule