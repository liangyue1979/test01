always @() begin
    
end